`timescale 1ns/1ns


module f_module(//output
                output [31 : 0] FxL,

                //inputs
                input clk,
                input rst,
                input [31:0] in

);

reg [31:0] S [3:0][255:0];

/* 
Check the python script.py for the S filling
integer pi_digits [255:0] = {
    3,1,4,1,5,9,2,6,5,3,5,8,9,7,9,3,
    2,3,8,4,6,2,6,4,3,3,8,3,2,7,9,5,
    0,2,8,8,4,1,9,7,1,6,9,3,9,9,3,7,
    5,1,0,5,8,2,0,9,7,4,9,4,4,5,9,2,
    3,0,7,8,1,6,4,0,6,2,8,6,2,0,8,9,
    9,8,6,2,8,0,3,4,8,2,5,3,4,2,1,1,
    7,0,6,7,9,8,2,1,4,8,0,8,6,5,1,3,
    2,8,2,3,0,6,6,4,7,0,9,3,8,4,4,6,
    0,9,5,5,0,5,8,2,2,3,1,7,2,5,3,5,
    9,4,0,8,1,2,8,4,8,1,1,1,7,4,5,0,
    2,8,4,1,0,2,7,0,1,9,3,8,5,2,1,1,
    0,5,5,5,9,6,4,4,6,2,2,9,4,8,9,5,
    4,9,3,0,3,8,1,9,6,4,4,2,8,8,1,0,
    9,7,5,6,6,5,9,3,3,4,4,6,1,2,8,4,
    7,5,6,4,8,2,3,3,7,8,6,7,8,3,1,6,
    5,2,7,1,2,0,1,9,0,9,1,4,5,6,4,8   
};
*/

initial begin
    S[0][0]=3; S[0][1]=1; S[0][2]=4; S[0][3]=1; S[0][4]=5; S[0][5]=9; S[0][6]=2; S[0][7]=6; S[0][8]=5; S[0][9]=3; S[0][10]=5;
    S[0][11]=8; S[0][12]=9; S[0][13]=7; S[0][14]=9; S[0][15]=3; S[0][16]=2; S[0][17]=3; S[0][18]=8; S[0][19]=4; S[0][20]=6;
    S[0][21]=2; S[0][22]=6; S[0][23]=4; S[0][24]=3; S[0][25]=3; S[0][26]=8; S[0][27]=3; S[0][28]=2; S[0][29]=7; S[0][30]=9;
    S[0][31]=5; S[0][32]=0; S[0][33]=2; S[0][34]=8; S[0][35]=8; S[0][36]=4; S[0][37]=1; S[0][38]=9; S[0][39]=7; S[0][40]=1;
    S[0][41]=6; S[0][42]=9; S[0][43]=3; S[0][44]=9; S[0][45]=9; S[0][46]=3; S[0][47]=7; S[0][48]=5; S[0][49]=1; S[0][50]=0;
    S[0][51]=5; S[0][52]=8; S[0][53]=2; S[0][54]=0; S[0][55]=9; S[0][56]=7; S[0][57]=4; S[0][58]=9; S[0][59]=4; S[0][60]=4;
    S[0][61]=5; S[0][62]=9; S[0][63]=2; S[0][64]=3; S[0][65]=0; S[0][66]=7; S[0][67]=8; S[0][68]=1; S[0][69]=6; S[0][70]=4;
    S[0][71]=0; S[0][72]=6; S[0][73]=2; S[0][74]=8; S[0][75]=6; S[0][76]=2; S[0][77]=0; S[0][78]=8; S[0][79]=9; S[0][80]=9;
    S[0][81]=8; S[0][82]=6; S[0][83]=2; S[0][84]=8; S[0][85]=0; S[0][86]=3; S[0][87]=4; S[0][88]=8; S[0][89]=2; S[0][90]=5;
    S[0][91]=3; S[0][92]=4; S[0][93]=2; S[0][94]=1; S[0][95]=1; S[0][96]=7; S[0][97]=0; S[0][98]=6; S[0][99]=7; S[0][100]=9;
    S[0][101]=8; S[0][102]=2; S[0][103]=1; S[0][104]=4; S[0][105]=8; S[0][106]=0; S[0][107]=8; S[0][108]=6; S[0][109]=5; S[0][110]=1;
    S[0][111]=3; S[0][112]=2; S[0][113]=8; S[0][114]=2; S[0][115]=3; S[0][116]=0; S[0][117]=6; S[0][118]=6; S[0][119]=4; S[0][120]=7;
    S[0][121]=0; S[0][122]=9; S[0][123]=3; S[0][124]=8; S[0][125]=4; S[0][126]=4; S[0][127]=6; S[0][128]=0; S[0][129]=9; S[0][130]=5;
    S[0][131]=5; S[0][132]=0; S[0][133]=5; S[0][134]=8; S[0][135]=2; S[0][136]=2; S[0][137]=3; S[0][138]=1; S[0][139]=7; S[0][140]=2;
    S[0][141]=5; S[0][142]=3; S[0][143]=5; S[0][144]=9; S[0][145]=4; S[0][146]=0; S[0][147]=8; S[0][148]=1; S[0][149]=2; S[0][150]=8;
    S[0][151]=4; S[0][152]=8; S[0][153]=1; S[0][154]=1; S[0][155]=1; S[0][156]=7; S[0][157]=4; S[0][158]=5; S[0][159]=0; S[0][160]=2;
    S[0][161]=8; S[0][162]=4; S[0][163]=1; S[0][164]=0; S[0][165]=2; S[0][166]=7; S[0][167]=0; S[0][168]=1; S[0][169]=9; S[0][170]=3;
    S[0][171]=8; S[0][172]=5; S[0][173]=2; S[0][174]=1; S[0][175]=1; S[0][176]=0; S[0][177]=5; S[0][178]=5; S[0][179]=5; S[0][180]=9;
    S[0][181]=6; S[0][182]=4; S[0][183]=4; S[0][184]=6; S[0][185]=2; S[0][186]=2; S[0][187]=9; S[0][188]=4; S[0][189]=8; S[0][190]=9;
    S[0][191]=5; S[0][192]=4; S[0][193]=9; S[0][194]=3; S[0][195]=0; S[0][196]=3; S[0][197]=8; S[0][198]=1; S[0][199]=9; S[0][200]=6;
    S[0][201]=4; S[0][202]=4; S[0][203]=2; S[0][204]=8; S[0][205]=8; S[0][206]=1; S[0][207]=0; S[0][208]=9; S[0][209]=7; S[0][210]=5;
    S[0][211]=6; S[0][212]=6; S[0][213]=5; S[0][214]=9; S[0][215]=3; S[0][216]=3; S[0][217]=4; S[0][218]=4; S[0][219]=6; S[0][220]=1;
    S[0][221]=2; S[0][222]=8; S[0][223]=4; S[0][224]=7; S[0][225]=5; S[0][226]=6; S[0][227]=4; S[0][228]=8; S[0][229]=2; S[0][230]=3;
    S[0][231]=3; S[0][232]=7; S[0][233]=8; S[0][234]=6; S[0][235]=7; S[0][236]=8; S[0][237]=3; S[0][238]=1; S[0][239]=6; S[0][240]=5;
    S[0][241]=2; S[0][242]=7; S[0][243]=1; S[0][244]=2; S[0][245]=0; S[0][246]=1; S[0][247]=9; S[0][248]=0; S[0][249]=9; S[0][250]=1;
    S[0][251]=4; S[0][252]=5; S[0][253]=6; S[0][254]=4; S[0][255]=8; S[1][0]=3; S[1][1]=1; S[1][2]=4; S[1][3]=1; S[1][4]=5; S[1][5]=9;
    S[1][6]=2; S[1][7]=6; S[1][8]=5; S[1][9]=3; S[1][10]=5;
    S[1][11]=8; S[1][12]=9; S[1][13]=7; S[1][14]=9; S[1][15]=3; S[1][16]=2; S[1][17]=3; S[1][18]=8; S[1][19]=4; S[1][20]=6;
    S[1][21]=2; S[1][22]=6; S[1][23]=4; S[1][24]=3; S[1][25]=3; S[1][26]=8; S[1][27]=3; S[1][28]=2; S[1][29]=7; S[1][30]=9;
    S[1][31]=5; S[1][32]=0; S[1][33]=2; S[1][34]=8; S[1][35]=8; S[1][36]=4; S[1][37]=1; S[1][38]=9; S[1][39]=7; S[1][40]=1;
    S[1][41]=6; S[1][42]=9; S[1][43]=3; S[1][44]=9; S[1][45]=9; S[1][46]=3; S[1][47]=7; S[1][48]=5; S[1][49]=1; S[1][50]=0;
    S[1][51]=5; S[1][52]=8; S[1][53]=2; S[1][54]=0; S[1][55]=9; S[1][56]=7; S[1][57]=4; S[1][58]=9; S[1][59]=4; S[1][60]=4;
    S[1][61]=5; S[1][62]=9; S[1][63]=2; S[1][64]=3; S[1][65]=0; S[1][66]=7; S[1][67]=8; S[1][68]=1; S[1][69]=6; S[1][70]=4;
    S[1][71]=0; S[1][72]=6; S[1][73]=2; S[1][74]=8; S[1][75]=6; S[1][76]=2; S[1][77]=0; S[1][78]=8; S[1][79]=9; S[1][80]=9;
    S[1][81]=8; S[1][82]=6; S[1][83]=2; S[1][84]=8; S[1][85]=0; S[1][86]=3; S[1][87]=4; S[1][88]=8; S[1][89]=2; S[1][90]=5;
    S[1][91]=3; S[1][92]=4; S[1][93]=2; S[1][94]=1; S[1][95]=1; S[1][96]=7; S[1][97]=0; S[1][98]=6; S[1][99]=7; S[1][100]=9;
    S[1][101]=8; S[1][102]=2; S[1][103]=1; S[1][104]=4; S[1][105]=8; S[1][106]=0; S[1][107]=8; S[1][108]=6; S[1][109]=5; S[1][110]=1;
    S[1][111]=3; S[1][112]=2; S[1][113]=8; S[1][114]=2; S[1][115]=3; S[1][116]=0; S[1][117]=6; S[1][118]=6; S[1][119]=4; S[1][120]=7;
    S[1][121]=0; S[1][122]=9; S[1][123]=3; S[1][124]=8; S[1][125]=4; S[1][126]=4; S[1][127]=6; S[1][128]=0; S[1][129]=9; S[1][130]=5;
    S[1][131]=5; S[1][132]=0; S[1][133]=5; S[1][134]=8; S[1][135]=2; S[1][136]=2; S[1][137]=3; S[1][138]=1; S[1][139]=7; S[1][140]=2;
    S[1][141]=5; S[1][142]=3; S[1][143]=5; S[1][144]=9; S[1][145]=4; S[1][146]=0; S[1][147]=8; S[1][148]=1; S[1][149]=2; S[1][150]=8;
    S[1][151]=4; S[1][152]=8; S[1][153]=1; S[1][154]=1; S[1][155]=1; S[1][156]=7; S[1][157]=4; S[1][158]=5; S[1][159]=0; S[1][160]=2;
    S[1][161]=8; S[1][162]=4; S[1][163]=1; S[1][164]=0; S[1][165]=2; S[1][166]=7; S[1][167]=0; S[1][168]=1; S[1][169]=9; S[1][170]=3;
    S[1][171]=8; S[1][172]=5; S[1][173]=2; S[1][174]=1; S[1][175]=1; S[1][176]=0; S[1][177]=5; S[1][178]=5; S[1][179]=5; S[1][180]=9;
    S[1][181]=6; S[1][182]=4; S[1][183]=4; S[1][184]=6; S[1][185]=2; S[1][186]=2; S[1][187]=9; S[1][188]=4; S[1][189]=8; S[1][190]=9;
    S[1][191]=5; S[1][192]=4; S[1][193]=9; S[1][194]=3; S[1][195]=0; S[1][196]=3; S[1][197]=8; S[1][198]=1; S[1][199]=9; S[1][200]=6;
    S[1][201]=4; S[1][202]=4; S[1][203]=2; S[1][204]=8; S[1][205]=8; S[1][206]=1; S[1][207]=0; S[1][208]=9; S[1][209]=7; S[1][210]=5;
    S[1][211]=6; S[1][212]=6; S[1][213]=5; S[1][214]=9; S[1][215]=3; S[1][216]=3; S[1][217]=4; S[1][218]=4; S[1][219]=6; S[1][220]=1;
    S[1][221]=2; S[1][222]=8; S[1][223]=4; S[1][224]=7; S[1][225]=5; S[1][226]=6; S[1][227]=4; S[1][228]=8; S[1][229]=2; S[1][230]=3;
    S[1][231]=3; S[1][232]=7; S[1][233]=8; S[1][234]=6; S[1][235]=7; S[1][236]=8; S[1][237]=3; S[1][238]=1; S[1][239]=6; S[1][240]=5;
    S[1][241]=2; S[1][242]=7; S[1][243]=1; S[1][244]=2; S[1][245]=0; S[1][246]=1; S[1][247]=9; S[1][248]=0; S[1][249]=9; S[1][250]=1;
    S[1][251]=4; S[1][252]=5; S[1][253]=6; S[1][254]=4; S[1][255]=8; S[2][0]=3; S[2][1]=1; S[2][2]=4; S[2][3]=1; S[2][4]=5;
    S[2][5]=9; S[2][6]=2; S[2][7]=6; S[2][8]=5; S[2][9]=3; S[2][10]=5; S[2][11]=8; S[2][12]=9; S[2][13]=7; S[2][14]=9;
    S[2][15]=3; S[2][16]=2; S[2][17]=3; S[2][18]=8; S[2][19]=4; S[2][20]=6; S[2][21]=2; S[2][22]=6; S[2][23]=4; S[2][24]=3;
    S[2][25]=3; S[2][26]=8; S[2][27]=3; S[2][28]=2; S[2][29]=7; S[2][30]=9; S[2][31]=5; S[2][32]=0; S[2][33]=2; S[2][34]=8;
    S[2][35]=8; S[2][36]=4; S[2][37]=1; S[2][38]=9; S[2][39]=7; S[2][40]=1; S[2][41]=6; S[2][42]=9; S[2][43]=3; S[2][44]=9;
    S[2][45]=9; S[2][46]=3; S[2][47]=7; S[2][48]=5; S[2][49]=1; S[2][50]=0; S[2][51]=5; S[2][52]=8; S[2][53]=2; S[2][54]=0;
    S[2][55]=9; S[2][56]=7; S[2][57]=4; S[2][58]=9; S[2][59]=4; S[2][60]=4; S[2][61]=5; S[2][62]=9; S[2][63]=2; S[2][64]=3;
    S[2][65]=0; S[2][66]=7; S[2][67]=8; S[2][68]=1; S[2][69]=6; S[2][70]=4; S[2][71]=0; S[2][72]=6; S[2][73]=2; S[2][74]=8;
    S[2][75]=6; S[2][76]=2; S[2][77]=0; S[2][78]=8; S[2][79]=9; S[2][80]=9; S[2][81]=8; S[2][82]=6; S[2][83]=2; S[2][84]=8;
    S[2][85]=0; S[2][86]=3; S[2][87]=4; S[2][88]=8; S[2][89]=2; S[2][90]=5; S[2][91]=3; S[2][92]=4; S[2][93]=2; S[2][94]=1;
    S[2][95]=1; S[2][96]=7; S[2][97]=0; S[2][98]=6; S[2][99]=7; S[2][100]=9; S[2][101]=8; S[2][102]=2; S[2][103]=1; S[2][104]=4;
    S[2][105]=8; S[2][106]=0; S[2][107]=8; S[2][108]=6; S[2][109]=5; S[2][110]=1; S[2][111]=3; S[2][112]=2; S[2][113]=8; S[2][114]=2;
    S[2][115]=3; S[2][116]=0; S[2][117]=6; S[2][118]=6; S[2][119]=4; S[2][120]=7; S[2][121]=0; S[2][122]=9; S[2][123]=3; S[2][124]=8;
    S[2][125]=4; S[2][126]=4; S[2][127]=6; S[2][128]=0; S[2][129]=9; S[2][130]=5; S[2][131]=5; S[2][132]=0; S[2][133]=5; S[2][134]=8;
    S[2][135]=2; S[2][136]=2; S[2][137]=3; S[2][138]=1; S[2][139]=7; S[2][140]=2; S[2][141]=5; S[2][142]=3; S[2][143]=5; S[2][144]=9;
    S[2][145]=4; S[2][146]=0; S[2][147]=8; S[2][148]=1; S[2][149]=2; S[2][150]=8; S[2][151]=4; S[2][152]=8; S[2][153]=1; S[2][154]=1;
    S[2][155]=1; S[2][156]=7; S[2][157]=4; S[2][158]=5; S[2][159]=0; S[2][160]=2; S[2][161]=8; S[2][162]=4; S[2][163]=1; S[2][164]=0;
    S[2][165]=2; S[2][166]=7; S[2][167]=0; S[2][168]=1; S[2][169]=9; S[2][170]=3; S[2][171]=8; S[2][172]=5; S[2][173]=2; S[2][174]=1;
    S[2][175]=1; S[2][176]=0; S[2][177]=5; S[2][178]=5; S[2][179]=5; S[2][180]=9; S[2][181]=6; S[2][182]=4; S[2][183]=4; S[2][184]=6;
    S[2][185]=2; S[2][186]=2; S[2][187]=9; S[2][188]=4; S[2][189]=8; S[2][190]=9; S[2][191]=5; S[2][192]=4; S[2][193]=9; S[2][194]=3;
    S[2][195]=0; S[2][196]=3; S[2][197]=8; S[2][198]=1; S[2][199]=9; S[2][200]=6; S[2][201]=4; S[2][202]=4; S[2][203]=2; S[2][204]=8;
    S[2][205]=8; S[2][206]=1; S[2][207]=0; S[2][208]=9; S[2][209]=7; S[2][210]=5; S[2][211]=6; S[2][212]=6; S[2][213]=5; S[2][214]=9;
    S[2][215]=3; S[2][216]=3; S[2][217]=4; S[2][218]=4; S[2][219]=6; S[2][220]=1; S[2][221]=2; S[2][222]=8; S[2][223]=4; S[2][224]=7;
    S[2][225]=5; S[2][226]=6; S[2][227]=4; S[2][228]=8; S[2][229]=2; S[2][230]=3; S[2][231]=3; S[2][232]=7; S[2][233]=8; S[2][234]=6;
    S[2][235]=7; S[2][236]=8; S[2][237]=3; S[2][238]=1; S[2][239]=6; S[2][240]=5; S[2][241]=2; S[2][242]=7; S[2][243]=1; S[2][244]=2;
    S[2][245]=0; S[2][246]=1; S[2][247]=9; S[2][248]=0; S[2][249]=9; S[2][250]=1; S[2][251]=4; S[2][252]=5; S[2][253]=6; S[2][254]=4;
    S[2][255]=8; S[3][0]=3; S[3][1]=1; S[3][2]=4; S[3][3]=1; S[3][4]=5; S[3][5]=9; S[3][6]=2; S[3][7]=6; S[3][8]=5;
    S[3][9]=3; S[3][10]=5; S[3][11]=8; S[3][12]=9; S[3][13]=7; S[3][14]=9; S[3][15]=3; S[3][16]=2; S[3][17]=3; S[3][18]=8;
    S[3][19]=4; S[3][20]=6; S[3][21]=2; S[3][22]=6; S[3][23]=4; S[3][24]=3; S[3][25]=3; S[3][26]=8; S[3][27]=3; S[3][28]=2;
    S[3][29]=7; S[3][30]=9; S[3][31]=5; S[3][32]=0; S[3][33]=2; S[3][34]=8; S[3][35]=8; S[3][36]=4; S[3][37]=1; S[3][38]=9;
    S[3][39]=7; S[3][40]=1; S[3][41]=6; S[3][42]=9; S[3][43]=3; S[3][44]=9; S[3][45]=9; S[3][46]=3; S[3][47]=7; S[3][48]=5;
    S[3][49]=1; S[3][50]=0; S[3][51]=5; S[3][52]=8; S[3][53]=2; S[3][54]=0; S[3][55]=9; S[3][56]=7; S[3][57]=4; S[3][58]=9;
    S[3][59]=4; S[3][60]=4; S[3][61]=5; S[3][62]=9; S[3][63]=2; S[3][64]=3; S[3][65]=0; S[3][66]=7; S[3][67]=8; S[3][68]=1;
    S[3][69]=6; S[3][70]=4; S[3][71]=0; S[3][72]=6; S[3][73]=2; S[3][74]=8; S[3][75]=6; S[3][76]=2; S[3][77]=0; S[3][78]=8;
    S[3][79]=9; S[3][80]=9; S[3][81]=8; S[3][82]=6; S[3][83]=2; S[3][84]=8; S[3][85]=0; S[3][86]=3; S[3][87]=4; S[3][88]=8;
    S[3][89]=2; S[3][90]=5; S[3][91]=3; S[3][92]=4; S[3][93]=2; S[3][94]=1; S[3][95]=1; S[3][96]=7; S[3][97]=0; S[3][98]=6;
    S[3][99]=7; S[3][100]=9; S[3][101]=8; S[3][102]=2; S[3][103]=1; S[3][104]=4; S[3][105]=8; S[3][106]=0; S[3][107]=8; S[3][108]=6;
    S[3][109]=5; S[3][110]=1; S[3][111]=3; S[3][112]=2; S[3][113]=8; S[3][114]=2; S[3][115]=3; S[3][116]=0; S[3][117]=6; S[3][118]=6;
    S[3][119]=4; S[3][120]=7; S[3][121]=0; S[3][122]=9; S[3][123]=3; S[3][124]=8; S[3][125]=4; S[3][126]=4; S[3][127]=6; S[3][128]=0;
    S[3][129]=9; S[3][130]=5; S[3][131]=5; S[3][132]=0; S[3][133]=5; S[3][134]=8; S[3][135]=2; S[3][136]=2; S[3][137]=3; S[3][138]=1;
    S[3][139]=7; S[3][140]=2; S[3][141]=5; S[3][142]=3; S[3][143]=5; S[3][144]=9; S[3][145]=4; S[3][146]=0; S[3][147]=8; S[3][148]=1;
    S[3][149]=2; S[3][150]=8; S[3][151]=4; S[3][152]=8; S[3][153]=1; S[3][154]=1; S[3][155]=1; S[3][156]=7; S[3][157]=4; S[3][158]=5;
    S[3][159]=0; S[3][160]=2; S[3][161]=8; S[3][162]=4; S[3][163]=1; S[3][164]=0; S[3][165]=2; S[3][166]=7; S[3][167]=0; S[3][168]=1;
    S[3][169]=9; S[3][170]=3; S[3][171]=8; S[3][172]=5; S[3][173]=2; S[3][174]=1; S[3][175]=1; S[3][176]=0; S[3][177]=5; S[3][178]=5;
    S[3][179]=5; S[3][180]=9; S[3][181]=6; S[3][182]=4; S[3][183]=4; S[3][184]=6; S[3][185]=2; S[3][186]=2; S[3][187]=9; S[3][188]=4;
    S[3][189]=8; S[3][190]=9; S[3][191]=5; S[3][192]=4; S[3][193]=9; S[3][194]=3; S[3][195]=0; S[3][196]=3; S[3][197]=8; S[3][198]=1;
    S[3][199]=9; S[3][200]=6; S[3][201]=4; S[3][202]=4; S[3][203]=2; S[3][204]=8; S[3][205]=8; S[3][206]=1; S[3][207]=0; S[3][208]=9;
    S[3][209]=7; S[3][210]=5; S[3][211]=6; S[3][212]=6; S[3][213]=5; S[3][214]=9; S[3][215]=3; S[3][216]=3; S[3][217]=4; S[3][218]=4;
    S[3][219]=6; S[3][220]=1; S[3][221]=2; S[3][222]=8; S[3][223]=4; S[3][224]=7; S[3][225]=5; S[3][226]=6; S[3][227]=4; S[3][228]=8;
    S[3][229]=2; S[3][230]=3; S[3][231]=3; S[3][232]=7; S[3][233]=8; S[3][234]=6; S[3][235]=7; S[3][236]=8; S[3][237]=3; S[3][238]=1;
    S[3][239]=6; S[3][240]=5; S[3][241]=2; S[3][242]=7; S[3][243]=1; S[3][244]=2; S[3][245]=0; S[3][246]=1; S[3][247]=9; S[3][248]=0;
    S[3][249]=9; S[3][250]=1; S[3][251]=4; S[3][252]=5; S[3][253]=6; S[3][254]=4; S[3][255]=8;
end

reg [31:0] tempAdd1,tempAdd2;
reg[31:0] tempXor;
reg [31:0] out;

always@(posedge clk or negedge rst)begin
    if(!rst)begin
        out <= 32'h0;
        tempAdd1 <= 32'h0;
        tempAdd2 <= 32'h0;
    end
    else begin
        tempAdd1 <= S[0][in[31:23]] + S[1][in[23:15]];
        tempXor <= tempAdd1 ^ S[2][in[15:7]];
        tempAdd2 <= tempXor + S[3][in[7:0]];
        out <= tempAdd2;
    end
end


assign FxL = out;

endmodule